magic
tech sky130A
magscale 1 2
timestamp 1756376748
<< obsli1 >>
rect 1104 2159 7084 8177
<< obsm1 >>
rect 14 2128 7806 8208
<< metal2 >>
rect 18 9617 74 10417
rect 2594 9617 2650 10417
rect 5170 9617 5226 10417
rect 7746 9617 7802 10417
rect 18 0 74 800
rect 2594 0 2650 800
rect 5170 0 5226 800
rect 7746 0 7802 800
<< obsm2 >>
rect 130 9561 2538 9617
rect 2706 9561 5114 9617
rect 5282 9561 7690 9617
rect 20 856 7800 9561
rect 130 800 2538 856
rect 2706 800 5114 856
rect 5282 800 7690 856
<< metal3 >>
rect 0 8168 800 8288
rect 7473 7488 8273 7608
rect 0 5448 800 5568
rect 7473 4768 8273 4888
rect 0 2728 800 2848
rect 7473 2048 8273 2168
<< obsm3 >>
rect 880 8088 7473 8261
rect 800 7688 7473 8088
rect 800 7408 7393 7688
rect 800 5648 7473 7408
rect 880 5368 7473 5648
rect 800 4968 7473 5368
rect 800 4688 7393 4968
rect 800 2928 7473 4688
rect 880 2648 7473 2928
rect 800 2248 7473 2648
rect 800 2075 7393 2248
<< metal4 >>
rect 1691 2128 2011 8208
rect 2351 2128 2671 8228
rect 3186 2128 3506 8208
rect 3846 2128 4166 8228
rect 4681 2128 5001 8208
rect 5341 2128 5661 8228
rect 6176 2128 6496 8208
rect 6836 2128 7156 8228
<< metal5 >>
rect 1056 7908 7156 8228
rect 1056 7248 7132 7568
rect 1056 6413 7156 6733
rect 1056 5753 7132 6073
rect 1056 4918 7156 5238
rect 1056 4258 7132 4578
rect 1056 3423 7156 3743
rect 1056 2763 7132 3083
<< labels >>
rlabel metal2 s 2594 0 2650 800 6 A[0]
port 1 nsew signal input
rlabel metal3 s 7473 7488 8273 7608 6 A[1]
port 2 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 A[2]
port 3 nsew signal input
rlabel metal3 s 0 2728 800 2848 6 A[3]
port 4 nsew signal input
rlabel metal3 s 0 5448 800 5568 6 B[0]
port 5 nsew signal input
rlabel metal2 s 18 0 74 800 6 B[1]
port 6 nsew signal input
rlabel metal2 s 5170 9617 5226 10417 6 B[2]
port 7 nsew signal input
rlabel metal3 s 7473 2048 8273 2168 6 B[3]
port 8 nsew signal input
rlabel metal2 s 2594 9617 2650 10417 6 Cin
port 9 nsew signal input
rlabel metal2 s 7746 9617 7802 10417 6 Cout
port 10 nsew signal output
rlabel metal2 s 5170 0 5226 800 6 Sum[0]
port 11 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 Sum[1]
port 12 nsew signal output
rlabel metal2 s 18 9617 74 10417 6 Sum[2]
port 13 nsew signal output
rlabel metal3 s 7473 4768 8273 4888 6 Sum[3]
port 14 nsew signal output
rlabel metal4 s 2351 2128 2671 8228 6 VGND
port 15 nsew ground bidirectional
rlabel metal4 s 3846 2128 4166 8228 6 VGND
port 15 nsew ground bidirectional
rlabel metal4 s 5341 2128 5661 8228 6 VGND
port 15 nsew ground bidirectional
rlabel metal4 s 6836 2128 7156 8228 6 VGND
port 15 nsew ground bidirectional
rlabel metal5 s 1056 3423 7156 3743 6 VGND
port 15 nsew ground bidirectional
rlabel metal5 s 1056 4918 7156 5238 6 VGND
port 15 nsew ground bidirectional
rlabel metal5 s 1056 6413 7156 6733 6 VGND
port 15 nsew ground bidirectional
rlabel metal5 s 1056 7908 7156 8228 6 VGND
port 15 nsew ground bidirectional
rlabel metal4 s 1691 2128 2011 8208 6 VPWR
port 16 nsew power bidirectional
rlabel metal4 s 3186 2128 3506 8208 6 VPWR
port 16 nsew power bidirectional
rlabel metal4 s 4681 2128 5001 8208 6 VPWR
port 16 nsew power bidirectional
rlabel metal4 s 6176 2128 6496 8208 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1056 2763 7132 3083 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1056 4258 7132 4578 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1056 5753 7132 6073 6 VPWR
port 16 nsew power bidirectional
rlabel metal5 s 1056 7248 7132 7568 6 VPWR
port 16 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 8273 10417
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 197302
string GDS_FILE /openlane/designs/rca4/runs/RUN_2025.08.28_10.24.21/results/signoff/ripple_carry_adder_4bit.magic.gds
string GDS_START 79448
<< end >>

